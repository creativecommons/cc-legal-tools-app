<!DOCTYPE html PUBLIC "-//W3C//DTD XHTML+RDFa 1.0//EN" "http://www.w3.org/MarkUp/DTD/xhtml-rdfa-1.dtd">

<html xmlns="http://www.w3.org/1999/xhtml"
xmlns:cc="http://creativecommons.org/ns#"
xmlns:dc="http://purl.org/dc/elements/1.1/"
xmlns:dct="http://purl.org/dc/terms/"
xmlns:frbr="http://purl.org/vocab/frbr/core#" xml:lang="sv">

<head about="http://creativecommons.org/licenses/by-nd/4.0/">
  <meta name="viewport" content="width=device-width, initial-scale=1.0" />
  <meta http-equiv="Content-Type" content="application/xhtml+xml; charset=utf-8" />
  <title>

  Creative Commons &mdash; Erkännande-IngaBearbetningar 4.0 Internationell
  &mdash; CC BY-ND 4.0

  </title>

  <meta http-equiv="content-type" content="text/html;charset=utf-8" />



</head>

<body typeof="cc:License" about="http://creativecommons.org/licenses/by-nd/4.0/" class="license ltr">

  <!-- RDF code here for backwards compatibility.  Please use the
       license's RDFa instead. -->
  <!-- RDF Generation Not Implemented -->

  <div id="page" class="site">
    <div class="site-inner">
      <a class="skip-link screen-reader-text" href="#content">Hoppa över till innehåll</a>


<div class="site-header-wrapper">
  <header id="masthead" class="site-header sticky-nav-main" role="banner">
    <div class="site-header-main">
      <div class="site-branding">
        <a class="cc-site-logo-link" href="https://creativecommons.org/" rel="home">
          <img class="cc-site-logo" width="303" height="72" src="https://creativecommons.org/wp-content/themes/cc/images/cc.logo.white.svg">
        </a>
      </div>

      <button id="menu-toggle" class="menu-toggle"><i class="cc-icon-menu"></i> <span>Meny</span></button>

      <div id="site-header-menu" class="site-header-menu">
        <nav id="mobile-navigation" class="mobile-navigation" role="navigation" aria-label="Mobile Menu">
          <div class="menu-mobile-menu-container"><ul id="menu-mobile-menu" class="mobile-menu">
            <li id="menu-item-48798" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-48798"><a href="https://creativecommons.org/share-your-work/">Dela ditt arbete</a></li>
            <li id="menu-item-48799" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-48799"><a href="https://creativecommons.org/use-remix/">Använd &#038; remix</a></li>
            <li id="menu-item-48800" class="menu-item menu-item-type-post_type menu-item-object-page page_item page-item-7466 menu-item-48800"><a href="https://creativecommons.org/about/">What We do</a></li>
            <li id="menu-item-48801" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-48801"><a href="https://creativecommons.org/blog/">Blogg</a></li>
            <li id="menu-item-48802" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-48802"><a href="https://network.creativecommons.org/?ref=global-affiliate-network">Global Network</a></li>
            <li id="menu-item-48803" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-48803"><a href="https://creativecommons.org/use-remix/search-the-commons/">Sök i Commons</a></li>
          </ul></div>
        </nav><!-- .main-navigation -->

        <nav id="site-navigation" class="main-navigation" role="navigation" aria-label="Primary Menu">
          <div class="menu-primary-menu-container"><ul id="menu-primary-menu" class="primary-menu">
            <li id="menu-item-48791" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-48791"><a href="https://creativecommons.org/share-your-work/">Dela ditt arbete</a></li>
            <li id="menu-item-48792" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-48792"><a href="https://creativecommons.org/use-remix/">Använd &#038; remix</a></li>
            <li id="menu-item-48570" class="menu-item menu-item-type-post_type menu-item-object-page page_item page-item-7466 menu-item-48570"><a href="https://creativecommons.org/about/">What We do</a></li>
            <li id="menu-item-48793" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-48793"><a href="https://creativecommons.org/blog/">Blogg</a></li>
          </ul></div>
        </nav>

        <nav id="secondary-navigation" class="secondary-navigation" role="navigation" aria-label="Secondary Menu">
          <div class="menu-secondary-menu-container"><ul id="menu-secondary-menu" class="secondary-menu">
            <li id="menu-item-55890" class="menu-item menu-item-type-custom menu-item-object-custom menu-item-55890"><a href="https://search.creativecommons.org/">Search for CC images</a></li>
            <li id="menu-item-48804" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-48804"><a href="https://network.creativecommons.org/?ref=global-affiliate-network">Global Network</a></li>
            <li id="menu-item-56460" class="menu-item menu-item-type-custom menu-item-object-custom menu-item-56460"><a href="https://us.e-activist.com/page/6747/subscribe/1?ea.tracking.id=mailing-list-page">Newsletters</a></li>
            <li id="menu-item-52800" class="menu-item menu-item-type-custom menu-item-object-custom menu-item-52800"><a href="https://store.creativecommons.org/">Store</a></li>
            <li id="menu-item-48806" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-48806"><a href="https://creativecommons.org/about/contact/">Kontakt</a></li>
          </ul></div>
        </nav>

        <nav id="social-navigation" class="social-navigation" role="navigation" aria-label="Social Links Menu">
          <div class="menu-social-links-container"><ul id="menu-social-links" class="social-links-menu">
            <li id="menu-item-48807" class="menu-item menu-item-type-custom menu-item-object-custom menu-item-48807"><a href="https://www.facebook.com/creativecommons"><span class="screen-reader-text">Facebook</span></a></li>
            <li id="menu-item-48808" class="menu-item menu-item-type-custom menu-item-object-custom menu-item-48808"><a href="https://twitter.com/creativecommons"><span class="screen-reader-text">Twitter</span></a></li>
            <li id="menu-item-48809" class="menu-item menu-item-type-custom menu-item-object-custom menu-item-48809"><a href="mailto:info@creativecommons.org"><span class="screen-reader-text">E-post</span></a></li>
          </ul></div>
        </nav>

      </div>
    </div>

  </header>
</div>


      <div id="content" class="site-content">
        <aside id="header-below" class="widget-area">
          <section id="text-15" class="widget-1 widget-first widget-last widget-odd widget widget_text">
            <div class="textwidget">
              <div id="donation-bar-wrapper" class="donation-bar-wrapper">
                <div id="donation-bar-inner" class="donation-bar-inner">
                  <p class="donate-text">Hjälp oss bygga ett livfullt, globalt sammarbetande commons</p>
                  <div class="donate-action"><a href="https://us.netdonor.net/page/6650/donate/1?ea.tracking.id=deed-top" class="button donate arrow">Donera<span class="hide-on-mobile"> Nu</span></a></div>
                </div>
              </div>
            </div>
          </section>
        </aside>


<div id="language-selector-block" class="container">
  <div class="language-selector-inner">
    <span dir="ltr" style="text-align: left">
      Denna sida finns tillgänglig på följande språk:
    </span>

    <img class="language-icon" src="/static/images/language_icon_x2.png" alt="Languages" />

    <select>

    </select>

  </div>
</div>


        <div id="primary" class="content-area">
          <main id="main" class="site-main container" role="main">
            <div id="deed" class="row" dir="ltr" style="text-align: left">
              <div id="deed-head" class="row">
                <div class="print-only icon cc-logo-print">
                  <img alt="cc logo" src="/static/images/deed/cc-logo.jpg">
                </div>
                <div id="cc-link">
                  <a rel="dc:creator dct:creator" href="/">
                    <span property="dc:title dct:title">Creative Commons</span>
                  </a>
                </div>
                <h1><span>Creative Commons Licens Deed</span></h1>

                <div id="deed-license">
                  <h2>
                    <span class="cc-license-icons">
                      <span id="cc-logo" class="icon"><img alt="cc logo" src="/static/images/deed/cc_icon_white_x2.png"></span>




                    </span>


  <span class="cc-license-title" property="dc:title dct:title">Erkännande-IngaBearbetningar 4.0 Internationell</span>
  <span class="cc-license-identifier" property="dc:identifier dct:identifier">
    (CC BY-ND 4.0)
  </span>

                  </h2>
                </div>
              </div>

              <div id="deed-main" dir="ltr" style="text-align: left" class="row">
                <div id="legalcode-block">
                  <div id="deed-disclaimer">

                      <span class="summary">
                        Detta är en lättläst sammanfattning av (och inte en ersättning för) <a href="legalcode" class="fulltext">licensen</a>.
                      </span>


                    <span class="disclaimer">
                      <a href="#" id="disclaimer_popup" class="helpLink">Friskrivning</a>.
                    </span>
                  </div>
                </div>

                <div id="deed-main-content" class="row ">

  <div id="deed-rights"
       dir="ltr" style="text-align: left" class="row">




    <div class="col-sm-offset-2 col-sm-8">
      <h3 style="text-align: center" resource="http://creativecommons.org/ns#Reproduction"
          rel="cc:permits">Du har tillstånd att:</h3>
      <ul class="license-properties">
        <li class="license share"
          rel="cc:permits"
          resource="http://creativecommons.org/ns#Distribution">
        <strong>Dela</strong> &mdash; kopiera och vidaredistribuera materialet oavsett medium eller format
        </li>




          <li class="license commercial">
            för alla ändamål, även kommersiellt.
          </li>

        <li id="more-container"
            class="license-hidden">
          <span id="devnations-container" />
        </li>
      </ul>
      </div>




  </div>

  <div class="row">
    <ul id="license-freedoms-no-icons" style="text-align: center" class="col-sm-offset-2 col-sm-8">
      <li class="license">Licensgivaren kan inte återkalla dessa friheter så länge du följer licensvillkoren.</li>
    </ul>
  </div>

  <div class="row"><div class="col-md-offset-1 col-md-10"><hr /></div></div>

  <div id="deed-conditions" class="row">
    <h3 style="text-align: center">På följande villkor:</h3>

    <ul dir="ltr" style="text-align: left" class="license-properties col-md-offset-2 col-md-8">

      <li class="license by">
          <p>
            <strong>Erkännande</strong> &mdash; <span rel="cc:requires"
          resource="http://creativecommons.org/ns#Attribution">Du måste ge <a href="#" id="appropriate_credit_popup" class="helpLink">ett korrekt erkännande</a></span>, ange en hyperlänk till licensen, och <span rel="cc:requires" resource="http://creativecommons.org/ns#Notice"><a href="#" id="indicate_changes_popup" class="helpLink">ange om bearbetningar är gjorda </a></span>.  Du behöver göra så i enlighet med god sed, och inte på ett sätt som ger en bild av att licensgivaren stödjer dig eller ditt användande.
            <span id="by-more-container"></span>
          </p>

          <p id="work-attribution-container" style="display:none;">
            <strong>
              Erkänn detta arbete:
            </strong>
            <br/>
            <input id="work-attribution" value="" type="text"
                   readonly="readonly" onclick="this.select()"
                   onfocus="document.getElementById('work-attribution').select();"/>
            <input id="license-code" type="hidden"
                   value="CC BY-ND 4.0" />
            <input id="license-url" type="hidden"
                   value="http://creativecommons.org/licenses/by-nd/4.0/" />
            <a href="" id="attribution_help" class="helpLink">
              <img src="/static/images/information.png"
                   alt="Information" />
            </a>
          </p>
        </li>



      <li class="license nd">
          <p>
            <strong>IngaBearbetningar</strong> &mdash; Om du <a href="#" id="some_kinds_of_mods_popup" class="helpLink">remixar, transformerar, eller bygger vidare på</a> materialet, får du inte distribuera det modifierade materialet.
            <span id="nd-more-container"></span>
          </p>
      </li>



    </ul>
  </div>
  <div class="row">
    <ul id="deed-conditions-no-icons" class="col-md-offset-2 col-md-8">
      <li class="license">
        <strong>Inga ytterligare begränsningar</strong> &mdash; Du får inte tillämpa lagliga begränsningar eller <a href="#" id="technological_measures_popup" class="helpLink">teknologiska metoder</a> som juridiskt begränsar andra från att gör något som licensen tillåter.
      </li>
    </ul>
  </div>
  <div class="row"><div class="col-md-offset-1 col-md-10"><hr /></div></div>
  <div id="deed-understanding" class="row">
    <h3 style="text-align: center">
      Anmärkningar:
    </h3>
    <ul class="understanding license-properties col-md-offset-2 col-md-8">


      <li class="license">
        Du behöver inte följa licensvillkoren för de delar av materialet som finns i public domain eller där ditt användande är tillåtet av en tillämplig <a href="#" id="exception_or_limitation_popup" class="helpLink">undantag eller begränsning</a>.
      </li>
      <li class="license">
        Inga garantier ges. Licensen ger eller ger dig inte alla de nödvändiga villkoren för ditt tänkta användande av verket. Till exempel, andra rättigheter som <a href="#" id="publicity_privacy_or_moral_rights_popup" class="helpLink">publicitet, integritetslagstiftning, eller ideella rättigheter </a> kan begränsa hur du kan använda verket.
      </li>
    </ul>



  </div>
  <span id="referrer-metadata-container" />

                </div>
              </div>

              <div class="row" id="footer">
                <p class="learn-more-cc">



        <a href="http://wiki.creativecommons.org/FAQ">Lär dig mer</a> om CC-licensiering, eller <a id="get_this" href="/choose/results-one?license_code=by-nd&amp;amp;jurisdiction=&amp;amp;version=4.0&amp;amp;lang=sv">använd licensen</a> för ditt eget material.



                </p>
                <noscript>
                  <div id="deed-donate-footer">
                    <div class="footer-trigger">
                      <img src="/static/images/deed/cc_heart_x2.png" class="footer-logo" alt="" width="133" height="117" />
                      <div class="footer-trigger-content">
                        <p>Detta innehåll är fritt tillgängligt under enkla juridiska termer eftersom Creative Commons är en ideell förening som är beroende av donationer. Om du tycker om  detta innehåll, och tycker om att det är gratis för alla, då tycker vi att du ska fundera på att bidra med en donation till stöd för vårt arbete.</p>
                        <a href="https://us.netdonor.net/page/6650/donate/1?ea.tracking.id=license-footer"><button>Make a Donation</button></a>
                      </div>
                    </div>
                  </div>
                </noscript>

<div id="languages">
  <span dir="ltr" style="text-align: left">
    Denna sida finns tillgänglig på följande språk:
  </span>
  <br/>


</div>


              </div>



<div id="deed-donate-slide" style="display: none;">
  <div class="slide-trigger">
    <div class="slide-close"></div>
    <img src="/static/images/deed/logo-cc-heart-white.png" class="slide-logo" alt="" width="100" height="88" />
    <p class="desktop-only">Detta innehåll är fritt tillgängligt under enkla juridiska termer eftersom Creative Commons är en ideell förening som är beroende av donationer. Om du tycker om  detta innehåll, och tycker om att det är gratis för alla, då tycker vi att du ska fundera på att bidra med en donation till stöd för vårt arbete.</p>
    <p class="mobile-only">När du delar med dig så vinner alla.</p>
    <div class="donate-box">
      <div class="widget-inner">
        <div class="gform_wrapper" id="gform_wrapper_10">
          <form method="get" id="gform_10" action="https://us.netdonor.net/page/6650/donate/1" class="deed-donate-form">
            <div id="field_10_1" class="gfield field_sublabel_below field_description_below">
              <label class="gfield_label">Bidrag idag till Creative Commons</label>
              <div class="ginput_container ginput_container_radio">
                <ul class="gfield_radio" id="input_10_1">
                  <li class="gchoice_10_1_0">
                    <input name="transaction.donationAmt" type="radio" value="5" id="choice_10_1_0" tabindex="1">
                    <label for="choice_10_1_0" id="label_10_1_0">$5</label>
                  </li>
                  <li class="gchoice_10_1_1">
                    <input name="transaction.donationAmt" type="radio" value="15" checked="checked" id="choice_10_1_1" tabindex="2">
                    <label for="choice_10_1_1" id="label_10_1_1">$15</label>
                  </li>
                  <li class="gchoice_10_1_2">
                    <input name="transaction.donationAmt" type="radio" value="25" id="choice_10_1_2" tabindex="3">
                    <label for="choice_10_1_2" id="label_10_1_2">$25</label>
                  </li>
                  <li class="gchoice_10_1_3">
                    <input name="transaction.donationAmt" type="radio" value="50" id="choice_10_1_3" tabindex="4">
                    <label for="choice_10_1_3" id="label_10_1_3">$50</label>
                  </li>
                  <li class="gchoice_10_1_4">
                    <input name="transaction.donationAmt" type="radio" value="gf_other_choice" id="choice_10_1_4" tabindex="5" onfocus="$(this).next('input').focus();">
                    <input name="transaction.donationAmt.other" type="text" id="input_10_1_other" tabindex="5" style="max-width: 80%" placeholder="Summa" aria-label="Summa">
                  </li>
                </ul>

                <input type="hidden" name="type" value="One Time">
                <input type="hidden" name="ea.tracking.id" value="deed-overlay">

                <input type="submit" id="gform_submit_button_10" class="gform_button button" value="Donera nu!" tabindex="6">
              </div>
            </div>
          </form>
        </div>
      </div>
    </div>
  </div>
</div>

            </div>
          </main>
        </div>
      </div>



<div class="site-footer-wrapper">
  <footer id="colophon" class="site-footer sticky-nav-main" role="contentinfo">
    <div class="cc-footer">
      <div class="column cc-footer-main">
        <div class="cc-footer-logo">
          <a href="https://creativecommons.org/" class="custom-logo-link" rel="home" itemprop="url">
            <img width="980" height="240"
                src="/static/images/cc.logo_.white_.png"
                class="custom-logo" alt="cc.logo.white" itemprop="logo"
                srcset="/static/images/cc.logo_.white_.png %} 980w,
                /static/images/cc.logo_.white_-300x73.png 300w,
                /static/images/cc.logo_.white_-768x188.png 768w,
                /static/images/cc.logo_.white_-140x34.png 140w,
                /static/images/cc.logo_.white_-50x12.png 50w,
                /static/images/cc.logo_.white_-270x66.png 270w,
                /static/images/cc.logo_.white_-245x60.png 245w"
                sizes="(max-width: 709px) 85vw, (max-width: 909px) 67vw, (max-width: 1362px) 62vw, 840px" /></a>
        </div>

        <div class="cc-footer-links">
          <div class="menu-footer-links-container">
            <ul id="menu-footer-links" class="menu">
              <li id="menu-item-48794" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-48794"><a href="https://creativecommons.org/about/contact/">Kontakt</a></li>
              <li id="menu-item-48795" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-48795"><a href="https://creativecommons.org/privacy/">Integritet</a></li>
              <li id="menu-item-48796" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-48796"><a href="https://creativecommons.org/policies/">Policyer</a></li>
              <li id="menu-item-48797" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-48797"><a href="https://creativecommons.org/terms/">Villkor</a></li>
            </ul>
          </div>
        </div>
      </div>

      <div class="column cc-footer-contact">
        <h6><a href="https://creativecommons.org/about/contact">Vi blir jätteglada om du hör av dig!</a></h6>

        <address>
          Creative Commons<br />
          PO Box 1866, Mountain View, CA 94042
        </address>

        <ul>
          <li><a href="mailto:info@creativecommons.org" class="mail">info@creativecommons.org</a></li>
          <li><a href="https://creativecommons.org/faq">Vanliga frågor</a></li>
        </ul>
      </div>

      <div class="column cc-footer-license">
        <div class="license-icons">
          <a rel="license" href="https://creativecommons.org/licenses/by/4.0/" title="Creative Commons Attribution 4.0 International license">
            <i class="cc-icon-cc"></i>
            <i class="cc-icon-cc-by"></i>
          </a>
        </div>
        <aside>
          <div xmlns:cc="https://creativecommons.org/ns#" about="https://creativecommons.org">
            <p>Except where otherwise <a class="subfoot" href="https://creativecommons.org/policies#license">noted</a>, content on this site is licensed under a <a class="subfoot" href="https://creativecommons.org/licenses/by/4.0/" rel="license">Creative Commons Attribution 4.0 International license</a>. <a class="subfoot" href="https://creativecommons.org/website-icons" target="blank">Icons</a> by The Noun Project.</p>
          </div>
        </aside>
      </div>
    </div>
  </footer>
</div>

    </div>
  </div>

  <div id="help-panels" style="display: none">


      <div id="help_disclaimer_popup" class="help_panel">
        <div class="hd">Friskrivning</div>

          <div class="bd">
            <p>Denna sammanfattning uppmärksammar enbart vissa av de viktigaste inslagen och villkoren från den faktiska licensen. Den är inte en licens och har inget juridiskt värde. Du bör noggrant gå igenom alla villkor i den faktiska licensen innan du använder det licensierade materialet.</p>

            <p>Creative Commons är ingen advokatbyrå och tillhandahåller inga juridiska tjänster eller juridisk rådgivning. Distribution eller visning av, samt länkning till denna handling eller licensen som sammanfattas skapar ingen advokat-klient- eller annat förhållande.</p>
          </div>

      </div>


  <div id="help_attribution_help" class="help_panel">
    <div class="hd">
      Vad betyder "Erkänna detta verk"?
    </div>
    <div class="bd">
      <p>Sidan du kom från innehöll inbäddad licensmetadata, inklusive hur skaparen vill bli omnämnd vid återanvändning. Du kan använda HTML-koden här för att referera till verket. Då kommer även metadata att inkluderas på din sida så att andra också kan hitta ursprungsverket.</p>
    </div>
  </div>

  <div id="help_mediation_and_arbitration_popup" class="help_panel">
    <div class="bd">
      <p>De tillämpliga medlingsreglerna kommer att bestämmas utifrån de upphovsrättsliga begränsningar som publiceras med verket, eller om inga då ska beslut fattas vid krav om medling. Om inget annat finns angivet i Copyrights noteringarna som kopplas till verket, kommer UNCITRAL medlingsregler att används vid medlingsbeslut.</p>
      <p><a href="http://wiki.creativecommons.org/Intergovernmental_Organizations#What_should_I_know_before_I_use_a_work_licensed_under_the_IGO_3.0_ported_licenses.3F">
        Mer information</a>.</p>
    </div>
  </div>

  <div id="help_appropriate_credit_popup" class="help_panel">
    <div class="bd">
      <p>Om det anges, måste du ange namnet på upphovsmannen och skriva ut villkoren för upphovsmannen, licensen, friskrivningsklausul och länka till verket. CC licenser före version 4.0 kräver också att du anger titeln på verket om det anges, och kan ha andra små skillnader </p>
      <p><a href="http://wiki.creativecommons.org/License_Versions#Detailed_attribution_comparison_chart">
        Mer information</a>.</p>
    </div>
  </div>

  <div id="help_indicate_changes_popup" class="help_panel">
    <div class="bd">
      <p>I 4.0, måste du indikera om du har modifierat materialet samt behålla indikeringar på tidigare modifieringar. I 3.0 och tidigare licensversioner krävs indikering av ändringar endast om du skapar en bearbetning.</p>
      <p><a href="http://wiki.creativecommons.org/Best_practices_for_attribution#This_is_a_good_attribution_for_material_you_modified_slightly">
        Märkningsguide</a>.</p>
      <p><a href="http://wiki.creativecommons.org/License_Versions#Modifications_and_adaptations_must_be_marked_as_such ">
        Mer information</a>.</p>
    </div>
  </div>

  <div id="help_same_license_popup" class="help_panel">
    <div class="bd">
      <p>Du kan även använd en licens som listas som likvärdig på <a href="https://creativecommons.org/compatiblelicenses">https://creativecommons.org/compatiblelicenses</a></p>
      <p><a href="http://wiki.creativecommons.org/FAQ#If_I_derive_or_adapt_material_offered_under_a_Creative_Commons_license.2C_which_CC_license.28s.29_can_I_use.3F">
        Mer information</a>.</p>
    </div>
  </div>

  <div id="help_commercial_purposes_popup" class="help_panel">
    <div class="bd">
      <p>En kommersiell användning är en som främst är avsedd för kommersiell nytta eller monetär ersättning.  </p>
      <p><a href="http://wiki.creativecommons.org/Frequently_Asked_Questions#Does_my_use_violate_the_NonCommercial_clause_of_the_licenses.3F">
        Mer information</a>.</p>
    </div>
  </div>

  <div id="help_some_kinds_of_mods_popup" class="help_panel">
    <div class="bd">
      <p>Att enbart ändra formatet skapar aldrig en bearbetning.</p>
      <p><a href="http://wiki.creativecommons.org/Frequently_Asked_Questions#When_is_my_use_considered_an_adaptation.3F">
        Mer information</a>.</p>
    </div>
  </div>

  <div id="help_technological_measures_popup" class="help_panel">
    <div class="bd">
      <p>Licensen förbjuder applikationer av effektiva teknologiska medel definierad med hänvisning till Artikel 11 i WIPO Copyright Treaty, WIPOs Upphovsrättsfördrag.</p>
      <p><a href="http://wiki.creativecommons.org/License_Versions#Application_of_effective_technological_measures_by_users_of_CC-licensed_works_prohibited">
        Mer information</a>.</p>
    </div>
  </div>

  <div id="help_exception_or_limitation_popup" class="help_panel">
    <div class="bd">
      <p>Rätten att använda verket enligt de undantag och begränsningar som finns i lagstiftningen, t.ex citaträtten, begränsas inte av CC licenserna. </p>
      <p><a href="http://wiki.creativecommons.org/Frequently_Asked_Questions#Do_Creative_Commons_licenses_affect_exceptions_and_limitations_to_copyright.2C_such_as_fair_dealing_and_fair_use.3F">
        Mer information</a>.</p>
    </div>
  </div>

  <div id="help_publicity_privacy_or_moral_rights_popup" class="help_panel">
    <div class="bd">
      <p>Du behöver få ytterligare tillstånd innan du använder materialet som du tänkt dig. </p>
      <p><a href="http://wiki.creativecommons.org/Considerations_for_licensors_and_licensees">
        Mer information</a>.</p>
    </div>
  </div>

  </div>

  /* <![CDATA[ */
  var screenReaderText = {"expand":"visa undermeny","collapse":"dölj undermeny"};
  /* ]]> */

</body>
</html>
